
`include "SquashCommon.v"

// The module in charge of the game logic, independently of the
// visual rendering aspects.
module SquashCore (
    // Add input and output ports here.
);

// Add module body.

endmodule
