
`include "SquashCommon.v"

// Define the visual rendering of the game objects and drive the VGA port.
module SquashDisplay (
    // Add input and output ports here.
);

// Add module body.

endmodule
